`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
bA3/TDYYAvcqhJsSQRf3H/hFBJMQlVKh1jhszAXMM28USs1PXlTeCqpfG2x+hD5iAufN91YD17zO
Bew+VgMHrllZ9JX8X49pqAmQYjl7fE/BUn+HNXHtst2NsL2nJpyZM1XedxIHmmlo+2QeHpDBRmeR
tVQCO1X3gq9vinmYdDdvzRsCn+lk848VBDAizJ5ru/J74IiAHmNN+ypt/o/gG7FSHWlYg6l20+T7
XuN4jTM7O4O36CYzAvvt2AvnsfgZaCrREg9LfUZMYy0gQBVRJH8TgkqzA6LrBJWn8uUmTFwESPoj
lsRmE0eXmlpNVy3c4WQQ4bOo6S84bFGPui8Ucw==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
VJYEGA6oowzFweH0iWgc2QSGRarY/gsU+hStDLdFcq/0TnsedTaoGeygLoJRsy1uCHXi/DC6rADk
EW3c79VodPYdh9l6Xy/9nO4UKseibPVWWq9245XF4iyTmvWymKXouuFGZvvsvATH6HyOTP9bhPAg
LCTUoEfjiIjX8qZhUh11kFuIR98VUODTa/V6/A1s1i0eVj4vzMdnmTM3YQ2MEEd7sgS9Di3OOCCr
51w2Mc4GjUoHEZzNshuuRV7Agsd9eNk4JVgadmWrxPkSmGthamn9AnL9Rkd+iQ04vzn8mJE/Je3s
RPtFLH2wlCtUhgtq/4Ev4EU19JXAeuG3vDL3QgAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FL+3W50R2W9SkvoqIXXv3vUO9dw+K8gfD6t6QCT+7F8eu8jOzIllKNx+uHAyeeU73iwxcKFlHnqr
6Nae4XgJAg==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J9dCY4ez7cwoor1/8c43HTnzjgqDzNvRRspyhpA0YIXFHomfkugvNdcqm0wEvjRFDqOQ32P02sWJ
LwoRDjcckuB3I10EuaDsLs9TFPdtr+pNjXlIQfW59cDhqXDQJDQq3t+9nZoDXrUvTRmQeRRdArRk
I7K5rjBatBIZG0j7Cw9+0Eo3AsUSXy2C41dG7tch7pdr/wA8xUf2Hve2QStABzK6F62BQ1iFpMZr
7w4r1zOr9DJX5d8QvVwfIU1u2+t2GgL2mkF66V9De+tr8I08Ztk7Z5K8q9l5plZ+wkgBSPs7pRaW
sl9HZ9L7MhzkkMGyMGjYru7OtMv4SDNDTIct5A==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
jurekguQgDQPTT2mx987nEjpKOSgr7vF6zfuq3ssrNuOd0/999JfJH/ETbddLBaXcOYvSITDlVdn
6iFM50ILw6qpbQ6tB6KRtq0qu+hinMnYlu321m7PzGDQpDK5da/eQCn0g37xgQwDY7kvvMpYQKLw
eOfdVzeP+ML1RMdVvaNNWYF9wjUaD8kFDXk7XQzNdRUGomXjzDzfe5FxKb+b8MqMyDo1kqYKRRq2
XW2Jk99/eRv/WpLy9x2wi+M1Xdjuxf6dfAzhLoM4QN92r4CeeUFEjnW/RomQ5nhxZCyPVI6tHLkv
HY3swWW7R2kmJNJBFpzTEJ6xVKXmOvNvKvbrkA==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
BknI/ebWkh8oDJa1F06uMO+iK+C3UpyrKGe39RVis/ZieJAIwY7vHpWbfONKcVwkw7YJFOAehYD7
amElWa2epnGLa+6HOlB/yZEZam2RpB2Fs+Th/JY2HOSAqcS0gZsesfEO46c7bOtccu77OyyBdMBw
/KTLDqtYZkjTZJm92Us=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
qVAWFicbcMbMKCKurNi1KGRzrmxO1PrmKQWQmT4rwsRbZ1Y8C7AL75nf+4ov5nIoLUY6L7qKdLjY
n1xRxlZlfJN80SEYncW9VG00ZaIPrPwsEKsdldz6wayFkXHfD+s5eGqPRjWe2a7Rq2h9hEvJf9CA
loX3YPfGwR+llUAAXo4KwyPXGjWTPHlXZ2CDA4r8ntr7L7XqU93+tWWovntDJdta4KHH6HH4wqHv
Cb0Qqr7tOVJ0YgICVVzNNXfvDkll+z1degXgzhnd7/4hmeXSy2OKjNk8MT8nJ+V39E43U1IefODq
+80TVwyLkHHRdoDDKdffjrT/tdkTZGrZ3y1Ong==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LXx2x+5G0KI5IEzOs653Si/YYcqULwUX1rMB+ZU+6gmFw6TrarTtKBP1JpJamTh1qBVG/OictX32
z3SPKaYwNFNzyLh7GC7Dj9hy7QDf/TkK4uRVmHm7goaTQBLP10mhp3FPPizXg7O0gg19JohYJaO/
iSBTRjAQE1H2UEMegbC8z9MDdBDakVrHQy6YJT/sUNsI3VzOiceFJOcWnBpP7Z0GFaGEumFrQ1ji
/FL1zmu7OfwWs8UaFZyyD1xfIoiFRsDN8CR+6ZIdEkUGBLq1d75Vr6M7re2GahUHz7j7eQBtFDQX
D3unf5/Okht1TpXi+FLQg6Rpjy5h9lYmNqSwxg==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
WrU+WsUptEt09hss47nGOjZ5EMMmJFh0qPj379Iuy1rlFEG6uPgaNdUC1Eb+9ILx1FHbqMwaI3MV
ZmrOEdO4emm0+0R/Dd4Af1CIHhwgcG2Rnf9+dBs8hJcFwLudJDF+1bnbs0ENP/U8Pl0jtTGkqdtq
+D2J8iSt8j3RDjf8p1c=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RNRa3/pBZdnmGjcpO0oNHqHXZX5BxU3L16+ys8VSxa1I3N8NOp8lSI9SbzGgbEQK1QhwTJ2cSeGE
394HXo+mEjddUpNB6dmfBoknMZvbXGiPyzxqfhua2RoE7puNp/EsfPL6qQF84at+qTcF0zSGlOhv
NFGVFa+3E9SoKmjNBUcqLtYZNkmhnnL/ZoWtOvYygTNdhaYNT/6MHL6wbDKKfMcEofUpSZFCEyZx
/HGbp9GeZjGuotqtgp/earZH9QVu9/9EYkJi9IPVwKpsHfohpCCzbd8ZCrj+7gfpFY/YfeXITs2C
dq7KKXcix3xTXIdWSngWzTNGshlTQuDR2sXdPg==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20640)
`pragma protect data_block
EtdDUSgARfq6GZOWeXZhSoDfV9A9gnSs8uPabasxHDsOnuV1iOC0WSb12ibBMP7Ela91JpXlugTC
h22hwwtB5649aoEYRrsgPOIJaHmrigPpsEgftUXGqQr3IRYhOhBQrueHfpo9No0XCCiFuNsoTOc0
IDB3rwNGYsXYjjFrxhPJ3rD5DA1lM+kIvoaHejn8FuhtABO5XStfRLWAvv5oTkN49BvXUGC+BmHr
vhqDDCmECCMS2g3M6GMpXs2EfKKAYS1rDUZAHyv/rRSuTW6RMdM7KxDIfQOUse1cnUSYoBusGc70
q5qKAORwMLtp3LMT30bfaBZeq0a70Z6wSGi58lbtzhEFybR5n8OBsYXTQCBfV6dCSvRH5yQouDwO
DgQRrltWwUJB+WxbAbrBDZp3n468L6nrptN0scqtZEN7JE2AZloWIr2jBfneFXY+Gm8JIq3kbRpU
3zahl1h1AVDolBAhrs5kpjw7JGL6TrcZBdgZHJqIYTd/5bdImj9UF93IFTUFhvBJ4xrQSH7u9mdN
8x3GQ72gZloTSMO2E5JYv528nFWztS9liBCwinPtTSJDpP4HhULBNDBfLhhzNPz3eg6K0r/iDVp7
PvM10/cAnTDRNl82OpkPtOnlh6KrqvMMilGAM/b0O/znHJ19lpWaO6C4de6TOUBIVB/Uc1/GKMo2
XrETeFdOQ3dUdVAMNJAIQ0cmjY/nvMRKrkdaSCBR5VrNYckOOo4dURWG0ZSQ6H1E4yKzNM3CLNM9
7gT2ve15v5SPjcpQsUjeWaA/Poztx8vWigp5UBx4wvxXhaMTt6+T8avEOtEaWMO3KpOYgpnQrwoY
a3ueTRxr87mBRYt8LhYGKaQmQudNnAZBwdzSSe7okquF5++i8pE5EM/6kOFY3epO4Q7SeNkw0rDi
rkBZNR7uWOBIYoRU88UKq3FPU5DIKy1y6DrNHr1WBVK6ZStpMcDZgp9h/M9TVmlowD1GZ4ZRutHp
y00Oubd2jYRLJo14IbfkBSEHFlO/f2jKv9Ypr1ZFR1Jmhlt6/iH60frUQ1LuCMOf56H1bHVZi3zj
0FPN4mkuw5A+e4tx7eIzOsw2UsQ5YgwSvlsCiJqbFvGgBn1D4P6rV7uAyCaxKmymn0+pxu1GpKPW
eCagBy8RQ1e2dWFFPF2qQsBYr3krZ3ront1Kwb/fr2OO01tBk6/H++O33kxYoG1v3V1FpnNRM7MQ
kQdzQsuYgrMmLKduxEwhAWvsQ/7U/761MPaCuS0fpqHBNDfOTxF38NpkG/V753R+W40W6Y19y5xP
DDN7rgZDk/nKUuvNBP7bUmc5/yjOHCmnhJh83isdrhA4+k4UxHVWaQ3Wh7Exx/rZE54jerjyNLSB
L2zewTisQjm1WyD6McjaP3vwpUevGXdfMgGEFg1VyUUQLxit0L/IovZgs93NMT4yLDEXzdF5EdEz
ny8fVe4m6SHNkIfTxBDP2DpTIA7joXGbryAp781g6/rM5MH5baqKGVKiU9znR+a5CFWV2FC0fU6r
4VPmUFBRj2kcOvtG31pPiBXgk6t9j91kJyRQkXDRfwvvdb6/FG82cjyZeLBFGWmYtjZeokJVXZN1
J9HrAcs+vOoew2g7VuHD3JynPAeY17tW1CXwQaK5mdM3AXJqeHbpzfBn3ARjG2SGusMQ6S/1a+E8
O/wjNoiU4/zm7GIvQaQVa+sXqvLJmOKk9k6nsQRiBUmHERtAIRjDyJajSY5WN9toLUAXUBTt29/z
RcxQYl1LZ+elRkZSxNyiivzFmzVSYSZSYvEK4zAZG+TeJl05taPcrzNYUSumUKnYBfCVZjnbfA+F
4COIh1cBhS/QC8QVRypplK8+vumHFjjnlTLBFUijoMa0yQ1JzTkRdPbgXO+W5fiu+dh20iyt9Tfo
z5tquZOUvJtGN9TRzATnOjNRPIGjnj4Xv53pEDuA4YeHJQjXOWyeAZR9QufWDqGtmB2g7APSeA6v
2BgUiei+EM0pNQWrcsttjOKl4gguB9krvDfAhL3vueT0oUI8+s+BobUAseq9MZvPBU/UKS+RNmkL
vWpFKnlNRt6Em+7Dk2PcpVVjUjeKj0FCOOCNqzqChojiJLkTiVZoGlg3Wz3aSMIZKA3fQQNfYPRt
dOdwyRu/fRUncb9wHvkK0FtvqHw+cCwHM+1SOZydKX5AXOA/zoTov38eY7rqmLyGszsqUIydr7ER
RzV//QHDeVttFGLzq3fnMP9Lman12k5yqRRE7EvgBJLi5H5OpYATeH0je7MG0Vy/ewzmODgoLBKb
heLfzkkgWVwsmPAAir57qlLAfziHJ1ngxwmlpn5DJ7weWMAT7FN1kMtPyTHJgwRcUFYmHnrT7AmD
R14xH8RzcBsQDY+eAF/jZZ0o1xC1Lx5o8uPtB2GYnhwUy1cGKFlEZrI5oW6SoRlW96cU/XOd4P+w
4Qaa63oEAFNTWLQxF2gBvYX7Cg2CKGhyLbkQ3qxPPoR1brqyGoV9yfQUPq0z+LxCLfsxuAeDow3O
2obb8s3YKlyFoufcYze78yiJk38woVF8P8vzEtkp7zHA7JYrnu+LERckHdANB+tp6CU5C39rcX3M
aNgPEjgo0Ou70uP1i7qjd0nDQMsN8SXGaCDnfbb1uXp6LyPxaDtnSm7SYsG8gHMqvj4bzhXbB8mB
mSQGrI0oESlbefC7yhuBaGXG20ydP34Kb1tufYQ5LIXB4WV2Q8ZGJCZhFL+4/l1jjwVtwrCnvLJ1
8/Ckc2hFQ2/g7XCtyZERxUilZVSasWynTXibIIL+LYizgyu3r8HrfKXCelXTeomQ4Qi1U6g13eaV
1BnrFrzlbONQ0TxOwFoTAa+ZYa43FT1pYTKG751Jpt16Yrt38FfYNEvsDne5lt4sN0OsOPs8LqIh
nIx4X9vz7a2TFfoLv4Il2Qy7E/F3k4/MTrwWTzeDg5R4djUfBgCTBu4L2UXqi7Oy6tRE2LQ8ng4F
sKnLAJ7beWKY/+Sk+5z6E1V52sAF7xEE16Ia1dX9L0jiMrPM/vmZJXFk58B+lXJd3YevBXN000sP
CqcS/8DPFy0K3CZ/1rTuA3XVfQBcJ5OBWZFtuT+D1yGChga5DQCfDJePQBC++isE9jaSdfyprbq9
DVTRaL3XREYMurxiBCALFygyfIXHtLsMwcANtA/SwNMx+y2/heQkzmBDwZ/J2fGy6zrByFQJEsB4
9l8vSaNCALmYd+fiEMIKKgiabTj+wF4NQarQwBQQWaq+Ly0urMAMTU7LRK/BkcdyPjIdLuiJwkdu
Nz0244iGFA2Y7/HtsPQ8fotDM2mnsTOEbrdwFgWEL72OSR5hvXe0fm/9PjM2TJ82582Yxd0n/C5D
4zLeoI0GG27kT5M15w8pwhcdwdPSFMDaMtUwMwSG9WlvPXBUDkFiPw8D77GuFW6C6XgGeQKYBm+O
WCTC3rB9BiyLBPtMwrYsAO/ISt9Gi+3Z+DjYFKKsR4wVhzNmLhNE6cdyT9W5QkYf/GynqmKtDEZS
FYFhTSU0kdfhmzSDJD6PDM88v/xtbnM5hr6DJa24Nmz/x2VRK5Qca8nPPvcCmo2p9CKSCof7aWp6
QX6whZ2tduQU+39/v0fI4BFaUivjw9m0PnFd44+tZ4t2qW8af3ECneRo2DZbfG1PQDtjy2zMBYis
SW7NTBA3QS3Zy32ePnhKEmUMGH7e/MEEV6u2l3KA16pt4DZq1dSaWtw+1iDqumqLGokC8GVKOe1j
FM7Gq3ZiUv72VHy3TdBb7rPCIWxL2b2mnDIIjqX1C2l+HeB9Gyc/ZEPLkPF7gIzENcg7QUsqNdcZ
HqHl1A525SwXD+993rxZvVSRci45LMhrRPql3Aujw30C1ReLlipJlLALSKOP6CkGk6zxwOG/4/cC
/eiQ6zB575lJcJtuPKyBC2p/JukjRGd12wg/QRZzt+G427WcFaKWbxEESQd0gqzsUtvCZP7GMfl1
T2xd63goI/repSQxYPocYIP5Ch/Cyu962f3uO1NzZkl7POw2GBuDbpUuY6GqCEjRVwFdQ05j7AMg
C3w0apiYIFgI4XoNaSk7z5evFQXEg/Y60jIqHNG6+RMCIgktXAhsmZOFOiq1sSnl7TexEyZsdgHv
JX3cdehhwu3cY5RMdGSiVWa9nz9gLpnBb+hVH9I2v3Io1MM5FlaSYxpI7UyjgnId1LRtHqbgwwhC
WO9ENPoQDaAC3Yrl7fA/mif85w+oROzyrc4MRmShnwjdarCAx5AvLgdV7CTUfeQDxihfrdKfv4Wg
I+iAxz0OhsJwIQ+vEwtkcGlM1VLU6wHzXn5P+HNx53Ft41/966YWYl4OjpIoQRIqWon9Lw48LZfc
sgE/BiBws8dWTFICVggM/ZgJ42nBsrolFDN/3Msz0eqpWf4RtkI9xxfNvkxEO1JwNAz1BIvHZn/A
o/p5l56FOui7GDzBbMHbsfxfiQN6jJVHsc5mhBCBAviUQaawpdMV/+/qotKlnwuFoSSFpVOt0vkM
44FBkxTAMJWuh1shuphMCWZ9oNty4IKgrgIPeGDLb6BBkfd96gz0k4FVI02SDfz21qWs9jCnuPzF
9L6Hl7fPEsSUHeoYmn8frkoFZ70lwamiPHkP0mVD1T11Atd6UTyT+wOTXOh/jhQIp0lwyVuqjnhU
WWFHAvpSTrl94FiW3kBt92plB2qZzAhXaw6fN3EhMmoTuEZzS9q7FfUxb9RLpwXcvaY3OYTW0CQ4
hOQh+e3vIBKpN9qyIpgTM0Ik1zdPoBIEzWQgW7HwJxeRzUtsULFH1IweLUsg5ixcLurezheup3xh
4Ee3otoNnPvLrXAUxRKLjkA0foxsdWuiVw+zTZXwd7R1hBEhhVT0mOf1fMgTpUDjGsxDGKHIxKhp
yzXkQ0t/ssIY9Zk2qkA1P2KFWoyh4k/2lfFiiTT7QYNZroYq5mz6jyCSBUzdnKK3X3W3GWaADsi3
J5LshkRIadivC4crXfZrSMkUKYXyLvaQz/atdRu3GGO33Z5xThAVMEOgG689hj+dKg7BQQXAYA0D
FA772PtQ836tM/x8ITvGQaBJtwYwxmugnbG+YhrJ6qwGpXDZ77hD22p4oQZfPwHTEFYU2BSTvOxM
vNb6jhifWPseB7FrEjlx80GA5eA+MJhfFIeonQEpwTC/JzFgG9V4/uCbzDIj3QF/sg8274Rr2Ieh
NQiilU+t0ppvWJ6Fczj/1PnAvbGTstz5U3rwQ0dYuH1DAz45lh0/GsoTfZlRD3PMB8AqEFkS+rYq
5ZhmwOCo00ihVy1S5pYwcfe4ECrXTRTvZyGQAduNqVuj8CEX/SIN4dUkSnOYRLltGy3jlSzQ9bys
vW3+xHb8IIv7vMWBDyA0rg4OvIcLPM8QUnl5ntpBINfhKOafwlX+Ba7jTf9xI5D09ftNF3LQtAac
+vbvyBsUp0ZAyDoU17d234c1c0nFDI4SWhdMqDsAR63qVmUihsLSU9Hq9jjQmLCeN2wPpcT0aZzh
YWgEn70vIpGS+cgCe4gYImpJ7cv94CDYADciuGNAMr8xGsqySPVpufpnexuqy3oPvRY+J6+xc4AH
V3X/oP7VwmN7bcac3bFhexP45qauCBNDG6prZPHYC5S/xFMSdvbhftEsR5gJ4GHCkFBozkEROtVg
JojzdKR5YVLI2flyB6JR6Ts7BN8gGaoA4PB0e9kxKPBD+W/5e7eVFCeoxQ8BomzvV5QaIHlH/gNo
CK9PVlqHvA4pfHjZfLCygXYSpHJhf+vnkZ933RmpR1YXGwpD69gYoYEGPal2IuCznuMBXioOG+5P
0m9a27BAT/6ddgbV10jdFiVsEWwU19+StRCRQBrXxD/YopIhpDSS8Qoi75YgggsxdxaBuPfiG1Nt
AOsdJ9FuP+kErTo3nxKse9ZP3ISQAoGLXQtoCMLdL/445Y9HNhyoY2JNs+S81LvknPbJY2kSCaUO
B7cPnXlWN0EK7+/YIZqtCJj0xxQS+LfIUSqXlgZh8W5xOIPy3ABXY7xRldh3uinunex8kFNjTmIW
dTxRK2MNAuvzL+WcJAnah6KWN3HPjlbGDKHEXugXLT40pm1P+6Cc1QhjdJOsT4Y1U/gk4xkOU1By
6BPmI5WxK0IKkOS/AFWl5v6ZA0UjpQlZ2LB11scqcf1gQ7q9PoqzBvf+7ZEJp8d9++osrTuDa84C
n/ouVFORe3ABMWy0ICZ84y3XGyRa6Mda+MF93BwmMJRmKWJHHmaa4u+yynCuWXrmVAKoZmoEwEXQ
RFl1KVNQeoj6Y20JDaHIXVwcPtUs46Asl6TZY2fxgl9ApbX5WtXQavPJ8WmBIPPaV+pyU34tLkQP
Ajx1RyjjJQtYpRRirMddrTk1RFLQxgxHVNxKRJoMyeYZtGCRQa2JJ6YLtL50/YD/pSVk6mwDyYrw
Lpndcz36Ne6Q7GOgr+tvGv6lmuCnJwBEXH+fnGETkJCScW4IWyDzm557R67dy/maDFrfMktqAS4K
YgaDqzspV2mqv2kNItfYmBDyoXIgzY+VGXWcoy3rV3fJ5/Z0aJDAComu9TjWKUbLZkPKNHkG8twU
nnzO9r4ArSQ7c/d++blAKZkf5qVa6yKw44NWb8WAojnH8iDym7U3LA3aAvUVUuV+PORIJ9jNPwv2
Dw3w7hIq6432hi5uNc/1BqODOGLsUAkKZ5MGlHQ667fwqE5q9USOriipXgIDYHJpvICv+i6F8xG1
UmFx+YFmoJHH9c8E4RJfJ7+UAASnXjUphJBQJOgW+r8CK2F0MLjWjsspGsVXsO9Z9G1ld5/Nrd62
srTR5CsWAfThjqrtVzZ7ekaDrfl2heYaSAAtJgSa8NiOA2oO85S79m9p9JcwaJC9TcG/+3fS4r/F
tcyMsKv0wqpI3pgn5/03nYVssyzdsD5daGALrXPpcyK7K8mM21Bngph072pRhjEDtpD7rHhgfDcZ
vdtAD4Cqe/EMx9h+Lje+5ozn5PIeYrgeLagp6jHjwMxM6NqBMhjC7gIDhh8OEnovHmSA7CqWHqkY
66rt/5YDh8ps9B9UkNZQzJyfpySSwOMRFZ3f/WRMt2Cy2K9BgQUzBt4Qgx5FfAvbqNQAdyhLVSFC
rktDKFHx7vCmXHK4okF5CH97qlhwPCdDK436+qLatSnZMWGU6IIEsMXF9V6+Ruqp782fPdGNUO7w
2nsbPSFEW5StOJR9z51QQ2SSZiFLGoeV6pWWj0tgoF9G2+CgVVdODDB8T4LxNnkmNhZ2vjjacRky
cSP8Rr2n0lltnylqHh6yCwqygg7uWgXFIlLFdoyyhQe6eiOV/KNFu0Y7XqyMoVAomfY+f5DpHllU
O5I5Dxa0XAFASM9nSr0Y0qTOfiCKCVbg7Af/0IC47DdH8YRhzcN4X0pFru5caiLEVutsK3SPYlQV
Iej/u7ViolZEwtuQyK3Puo3gYi7kZhzBqAv1xvkvAa/FBSL/X45vSKVtMM1sbdxFePUR9LA9s8wN
Tuj68YgTWZ9YM/xatOKqjXczsCKZQMj2BZ9rmrYfraO8yBm5VYWSpe6PZgd0jQ0NgwxAm3waJ+kL
LvgiOAL+GTowU1Ftcxf6n+Qe8p7TU8hcjWw0MxKyvwLUdXwQRAG6A/EWyrpWBMV33fMaWAmL4HQz
uZGeQJ9NhjHqDOzHPCq6GrAd+n3lJP4wn1QLD0CKbxj+zt64qGj+YLLxT5gP5sqfmGWHfPAT6YvD
OKXWANh6HDzbYs680MnOO1SzrgXwEneedYkCsm4/f9S5wIxk3JhAVp2QMpMdktMPtLe0iRToyXxC
p2blN61aaynLDgdj64UcHwA4DNuPIlz7SKwYdMrjWGSH5qv+sOhkA0KwgK7mY3UF6Rug916VfEC6
aPi8kWtft0nTOb+xIHDpCu4DCt5woehCd595mkJ3EIcN33xX08o9mX7PkH4jel/McNxPkYlgaVcN
C80DuzU0xrcPWF1eHvy2b7pVO7ZRe+KBPY58NdSoP/d/LO0qvA2cSLkpyZMMDoj9JSY7n1VsQ6qA
J/+eePwHug5K369q4oRIxMWKsbcWPehgBpmcaSO9ahcVcku7biz+LslWvCpV+Md3P/mkjGVMiBW2
J+XKAWKyTWHmHKODYLwC+APrXDJaWIqsRg5tk3jv6Xs0FJo25kqUNJbyrd38nTwjp1D+E/QbTG+9
NhDotBG3FpoqJuEhdwgmnBziS9OOntRVj1V9MPRKPwwbyGmCIYnnYZrJRUSdowC0JnnaIC81Yg2d
KE5doW+sPibFaBIqXiE2c9EOEvHyCes2VN4DWpa4nmXO0g9WhTsCL0YgdFbohcpxbEj5kPfo2s23
G8oy8j1D/kpexVdUW3VF+Y6xkWE9XPlV9LXD97hQnXKnjpYB/EPASLt5sEyxDOCsokGDvu8qaygG
k7NrHRtrZ0o5TLECdypUShY1XDHXR6dL8WcqR2I3VQR66+GszGz7qKsdiOgt8+pYOtIpSNlqh4zI
oFt8gP3psczaAVSntZ4ZY9kVQXYLYyMf+2efaNsPR9Rp9QFu8rAlP4yE+Oij/Y5PFqlRpfPMn7r8
W9NQFvDwsKP8awJayz2Pwec4DIyIvArJmQmI7x/mflIgwdxdjygRwMW9J+YMsP2Au17zcvjcuJEf
C/0D6aRDgXdIDQ72PN3AUw63mMWWY0Wol04RXvnNuKDRbuGKoXC8h4ZTZVlPFCTDzVLNXZ7z8X7d
BWUjlOJ7U1XyiTZ+Xqr3iS+nSx3IfOcJ6mbA4mVpj8gP+VZ7F20GwP+jlN+sfZo5t/HmLPVNQ1Ab
YwhIxmdmy2xrXPslfm4+mjjmhme7SmYMGSyaejVHOktSShkFW7j1K9HeKtYjJPMw3me2zPYGL3Fh
r4GN49dNKzzxWWI4KgrkBDfE5+6ZotzQAictbQfKJTbM0xdUVGtOAwaJut3sZKozzUAv+9sHwdrA
inao4IlYy55aiX5T9uSn+jjuRW8Ez40MsLd7/pX6de5vcvpGeZjY4yvqh+hiH5MybXGzb0GPDAXf
EDiUIzpnVRcyumo0iuRAPWXbWr7Ih1ecjKLN9h5aXS5GxBxfqWcxgPFkC+lum4D5vOpWy/Lt6YFl
INbFE1ARj8Gaj90vYejc6TO2AP89vgPjXeZi5ikSXkeZBh6rHYLH2/NTpZRuISzfe04R7pmagK9a
GhZqiFhTikpZrAVqekzeKytyHk2kEWGrlJZZlr1IikqOu47/WPsj+1ei/zEjIFwfmE8BoGh5Y0lM
PNec+SA3Rqz9JlH6wfBCGfqqFNFhJdn3/GljGFgYaAJwYFD2hEe+Wa5YkTmrEsnuTzMSrlqfmsL0
Q6vA7KlrdSRjYDXmHkbs/TSzhCTt5TQu3a9LG3IOsGboJupHX/BiK1VKc98wBMOinEB9j/92Kq7G
8xijfy4vOY0OJWH99TPrZuawSR2yNy+04w0GRLKjW+HaxN2VI1Omar6ncxeA5cgZYd1d/kU1BEZp
u8YynAENJxQp5ism30UuU8USZXHaQPLD0Yq3GmkdOSTY6B3tsC9SM3MQewNXisL58gp4GklAoqw1
CzQa5GJJ2T0+I8vKfP2UhVNbRRE8DXhzCsJ3exdu6AZfvzgEOOp11ZP6vbeYpCLenYvLl9+tOhwu
+yU8ciNtNCXMVhwyWrWQ9OoEB36yiXnfDnq6jafirkk7V5s3vB7gpCF6OdG7JeKuXxMKjbnWdOoI
Xk9BqMmQ7OAHHyUi5DkId/o3eUpGHQoED2tYJASLZfDXOLrjURkaUaJWd5MYFwAVJzixxy34kdpG
WfKjaZfb42RHrbSkeNaaLVjeIcv8bHb8hfshv9u6zA0fSIKl2pbkgm87bcjLX1AqAKcowGCb00uD
V9hCIwbVb7Ge5aKGCJafGHz6H9Vn9/kXEpB7qJCCtctQFQAdsNXBJLTxcdQ/oInS+rqrUPGL0YUx
ZLIAYp7AmiSwejpXwGRf8lvJdQoKyj8ehehZ1dY49WtiRxd0yIL2Ynqv9vQ3s9qq2KC4Fy8PLCYQ
wWlIKFW3eIqt4a68YOwhzs4TmV+KetizseD2XwWhWu50QEfHvGb0oVz8r5TrKqTysunGFX8GkXW1
A/qrLdAe8J3zljdTqNNUtexewRe1Nvnac9TDnT3pN2+iKsJyZJ2xEm0uFwoIW7+n7YMsdYKRqJF0
96dk9InsCujIkSFBukUt7LnSCHGGWoj4auZm5jKTSVWFoD1VmWF6sXpuqczPF03USGVGfz6S4ctz
vaty3LE5wdfKBaZtnJMvrH8f1rpbGneeeU9nHWfOuCtpEZJrp+D0usSkv3HeLOmXACxjxYCWRLbZ
QVjSLVF7xzDkmMfiTpuKigtDAQsnwS0vyjvkLxyOXzhjajgjeDL3OmmHvOtppyXtj4YKmnIaj+b3
rySNjCUds6JGF4L2gE+dkbbLh/AuVPUTskawGUW5AODcjhTSfjhw8NPo7hwyZfXSjFqbbC7RVB7+
OHe+p2g2HIjRzehl8twwAfKdKwKn5qYq1nvYiIOjK3UEXB4lLpVm+XBKDaBLrtvdYhFeAqJJ9SkS
b3d4jUxdEOT6Fl6SPcsw8G8W+7xvuXPg5fjKlEewjdWtXapHStIKD5hK9b4glcMb+1t0i4zWzE5I
/cPx4G6WqWdf8eIT+SAAw/f37CBnyhJNI5Q1pqgqfonD2ygPLeZqivL2StuJEmMvpJAnWcYt2047
NL4LHjOtx3VKPUeQOqhMyYKDnme4R82PZpL0/Pgp8Ra/rlaTt/1hClQ/6gVXuuFUP63GYQjyEcrB
VXzVmUvDede+/Dl8Po54YXmrXaXgDeR182ziEOVjgy2gfqJBtOxTgx89yZir10h+5hKE2DKv0UeT
ptFiT3vp1wFcvETp0NUtwlGA7fMTDiHzJITgAvAb5OJQ2197DQlGf6KXMlYGNFmzV8GHsMZfr3QN
gB7ID9GIXK9Md+slpl9QwfDpO4kWH6c1gQip7hnyikFWNECuhYz3owl2YC6WwB4vPmRJFrrutJ01
BBObsWDIK73sHiEXhtiGW+4tbSlBLxM6jYL2V3i0jDZEPcb2cMZPpFgRRRgjC7hNPznugKyiueFh
l//CavLro9AyYaZkM7qunERfeRI8MdRRcTHJTDWFYaVXMGghJr6NeKkw9QOXnrG9wxz2fWVIPW5x
3V4rXhlZBlHafRQCl3fA0QrkmiLfV3pdzGj+6MZJGH6sgC1iOv6tc0AeaZuWtE1RaDGH8+Pc06Rg
f4eFgCMKgYwqiJl3xBFdGHqWx3ndSAkP2XsxJ950hC+yxfjDTkDVX14ZqM29KkvgMBB5xW1TgEXL
JfbJl3bpv06XtSAhleII+cwf1eY/9Xf07075noy+Wsei8PtCOt1d8ZJN+aKDXzujNNawdigIuVrt
PmePsM4lX8hV1wJ7ZyTG9RJYnGr2/H8doBHhC6Xj6/xbcP3SZeJISj8m+4WREjfZaapKlCoJuDXw
yz27UkXPXeDo0V3HFFakHTrEHPLF0GPoY1H9XhL4WBFeXHWO4fBrx6/ZeHvhvvAP0/CpAZUxjox+
F6w7QuNp67w3MDxIyfwxN59cUn6iXF2/X/CR2iDrMb2OvU5GUw6zwN+MHnJGnAyGlEskwop8D+Mg
i6xF2J+s0o62RQcttvk+xK2lQqRXvKfD+n7dCtESr7EmJaF+8DLHdFrf1cGM5FeujahdUzz4mcz5
EC+15Qmd7Kz/+i8JLgzbzLHyeqmECVnlDEnaFZby97EvdcbD+s0OZ0jLYygvufhpUskF+qHgv1Fx
tvXejb7AeYUrxTuR6X9kVQmlnff+63nt+AyosHPcUgEWXJGU919p4oW7Oqz6+aOneRsyEKehH+Pm
oS04GTOYTWCZziBaDmr/WzaZSXjDrh5SdgRqIL6BlXwDOu5GqOjZYCKAtFHtg5z///dAsSxgINSK
lKZepRRNMUnBdjHvWFvrS6yLdxF8lZeW9qCniFOk/bIZEhVjKIvWp+Wzl9fGV1Dw6Lp+vdV4TKSh
isMx00lvYmD+xj60S1RwqiGjwJsygShAF8RA40L7C6duQG0A30CWAXsKJh8ba6XypG5ng4Al4hqY
VG69kxiZ+ENbDNpPcU9cR78HEkwOzVIpUSLcYmNafp0g9ec3uCcEi/pyla6qbX4t3RxGt4RKZal1
+KZhnNI7Hil5wEOQ2QPbHz54ANrtrkTtKohgSNXC8skw4iJiWhtImMwpK75Q+aPwWxZp4Rn63N1M
NgBlkh/1KR9lIb9MKtTPK/ceZIorfoHpl82I+J21kqfPKeDYk/6qlYDi/OjgjzbiknDjPwJx77Y1
vgaduD264LDMDqAhvyoXVa6jzfpLUPLB+FgZfQ4GRd6krQ7PCqBrhUF3DE1W3sLQi0A+XH0eh00U
rrlGJwHTtIyTPaqCuga3o/Z19j8ikwRppsY4qXEC654mCede+Dk/9zCLd12g3cWEGgjvN4s4/OuN
0hOGMGNVGftDIly3/XqezvuuoX7Eoc8wcwXOmhV7UsslFCC3chaxZ92BxG8jTduOLhof5tDJpu/W
ixfGvuIbyYNk1eaohfSMNRi84hXAbYIHE1GkFeHEkkQLKJxN1Fmbb9KWpi56taFGhcbHswfvDu/b
Pf5hC0ChI76895fflRCT6H/hYpV9KAc2t+KfwtaiYGSeE6mnBJiRBgUaXcnPVH6LymtjLLv+p8CF
jhq/I9LFrxmbO/JEpIV+gggft4YnPFjIhvKQrn6wCxUA5ppLVWDKIzprM1r9CaOTIRh7HURDCkMt
5bO4Xu9Fh6A9r39UDS5ZBJwbPR9INM0GSxyMpkVCsQOqb2/dTQQyPdnVr4on5xSVlsNv3VB6Rnju
tHixNNqZ+L+ZWaBKWPe2G26jgGbM8A5kdouM+9EwhZkH18z1adKBjGl3wRWgCwddza8hqoFgWs4d
c0O1HT6VTy3zf9mqbS1Tfk1EmOktO8qCdVxYgEai3ejAe658HtLmhXh/W6RzHQVRAg58YnToRHHc
kD9tOHhvd2GQLqEcGid3yTgwB7JJkDJ+MmcorjS75JIeCMarLwNtbJOJ0oxBw2YQT/i4kd476z2o
Tf1N8Kb0oX4g5BPQLB2ckmv+OQ2wBrK+6nTQg+QXc9HsN0R7DspdsAlYgmXqzhBKervzD4la3xeG
VZhfkZepeCk7tJN2p+IA+dTvt/RHLpah6E0R2PRcn5lvC6wtdf/ItrS9mNmMISuy4nNRkLbD2mnw
3lf/2miHg6qOStQPdAKHu/bqUUPahi+zcP+WYUR6LqxbHFiwE47tE9Ut/9pXpwYPxhjZaq1NR1c2
e8FJiVQHPCMLphxOrtTAt5Ho6TSrcjOFHOjIKeGBWPNLNcaKILnu9l3j0KWkHUi78BA8EEyyroqG
Okn3/JDCuzOfeAuM5dYR1Q3DiHIRXzBW7foLDX8nmK3w0iGVyeBHyuMsyNgE0cOg4SJk+hf6g4OA
efFzxA0wMEPi6bwsKth3/TGfzdTyQVgpHm7WMcNYCRiLh3NINdgLZhBAt4ByFBlsOrsXp8f3KGOD
kH1kSPq1dluqd7sTlm/MjMAH0t16ep5DwoV2LNODCLx6VBLkTbECE3oNenWalStcSdtaIM32Ek03
TqOpJLonv3my4cPu8Owvtwi36iNXHDVgueVGmlNNrnn/ZDFBLDwgscINzAeIJ43waVE0CH8troXA
nYRHfOsGDRxGmcHPHWcL/zf92cf6fua27ZvEIdZUZcWq2mGdkapNIP/q4VLNS+e3EFmqti+DTr45
38Qv4s9uLK9uCyZySM3qsL7YR4sfV6f1uj6MoTahBAi5Jloa4bO2vK8XYXCrEBRZE7d8yTtk/cL0
U23xTtk5AybxQiTEwSqxj6ByOEmipqqwCkpSE/UtEDHL+8t2QCDz416HVxJwj6bWE3pUIREhcv8i
gdF9o1R/2uuWP6zYJNXGDeR/MvHJQTN3JlIleOBcR4ehH00dxvZWHjSWpNtDuJ9/xstaEbawSDEv
UfPo/MwU2Y0XhJiRHvNK12ryf9c29lIuXyMqMR1dnvmYOHcwNCtwo5g9SHRTwv04mun8Fpf4kTjI
RmUDydKZ3sVxMDTo7o8NKeqrEGHtEx5yk38P2cvQe37T+O7B6/HTvxeU9FgcpM7sGfzQP70UGplD
0yELFmxdt+g4Pz1XpjSd/4zeVFdgx6kPWCf1Qhl2CKu9rYJO7SabpJMUcOHteNPlljzSNrg9AV97
NEIqm2GzhdENsS6Vm0jjbOxgfPBr+evxVhDXMJeaEB3k4ZlnNmVNHMQdSEBxra36I9weprDxV0At
uFXF2rIxJSer2vgq/KP7lZPrB/EqQlC31xZz37BcH2m5wj8uLGL1dFqez8QNLcCxanUdSWoYnOnB
nRHhSdUD23dSd/FIOCjVqaHyIaB834KKSf51BN+V6sKYge5kb6dmQHd5RtOewaEsXyuCyMOrGFLk
khgGGLzH4iQGU44j7AM08X22PiM5rAOkxP/iIJSZrNDkYyZn1zJQjhgoVxfTnRR+sC4KvBRyI6nk
FCq2+g+r9E2/5FgocKvymNuQAP10mZ2A10nGw8FvMlm3c99itBtJ/TL7p5zQbyurEvxmuorJQ3xm
NokXRdNnJTLAB4/LHOaGz83zjLWR3QiXHGQEP+NaVSMplsbjYc3RsjZj3axxCmHbHQzQlwPtQExL
lU0zq2nLp6jg5gqUYpDuVGwdFScxgNhk78xCraNAQBpD+IzCTqdP7BPP3NzW45Ig2eYSA0PsxXq9
dWRG3x7YjblVP376/baHfuaB630/II2sHJQul9WG4ayVwdHZbutdI9Rl20pxhdqGUZI/MP0D9z0j
oaIy63n2/LQNyuPSj2WsoIz7IgVsjOraxHnmHx4qn27AsbhtCu+mkWVEb8+EmErosoIt4/c2/9OG
6hYpyHJ4IMYElrGK+8BzRAiofZ/sN5eYVwBq+aGKbMudNU3veVjMlZ217CorTGihmIhGf9HK+4fg
6d7uUK2vseVd1a1vrY2Uk+pXYLUfgznJcu3W4kD1lLoYgwzrkC7KETbmpzCDauNFJnLyyv8XRE6B
64VNNCuTsvusjn74YOUunn8p3DSH+43p6alnEONH3pYiHqpOwzMWVX5txqDPikutu991Zrz0/6rh
B+svWPFgVIDvJbSXusTdFG+5peuJLmbBL/MJOxK8PMc8Spgik+YFhhrTX8KXc+sDIW0G1nttFjti
tqhbci+/soY65cqdVjUAUt/VBeKWYGhdXizi+Y1Cb/GUdT1MQ04lYYW8hwo5k6MAHnvBnapYfzLf
bqjBBofDTM9gY2jpVFRxnHJu7hisHKlXMgT6ngsMYewx66K0gnA/dSI+9aRBu+ZzQzDZ76Ma1fBQ
gV5lSYcikQevBdlLCx043kdkg/d+a1fLsd08F2OpOlxiZBOd9LYjDALjMdf0mIur5/HZD9qGgMII
Eb88ZQL2i2lTyz4fkty3EZKpshteDQBTM7gVVT2kMViuDDoVzf5+uYncY6kQ/K7TZyleP+U5Zjf1
Vm4g6iAh48/v4hKCag3zI0QLurWoD6VfHGWIyFW56zcHRyioymmPXCWLdRZTF2AmLlQQT9IZSD1w
2zFmzokvBnXNVsgYxz4TKS6cFY3vp1RqjNuONEJeWQobbdlDNHV8s3zi5b4P+DSTpR1VrawSxbjG
CZxWbG4xpBh3CnHWBiS8z8XnFbZzwCBwW7YKsNha5AIGjCXvR7CELgG6yRqFDucSDxSLkOfE5ih4
k8gF4s2g7jAKnK4sdtGQDwhp6upGAFFG2MNmW+59spwn/r5ahSE5ErtK+Bola8ncsbMuy8ZZxT0c
BbrZCWIGC3SJpamBrq8aMNSib435tc9uL3plXlVtqKj9PBWxb7jxksYA9bm9tXQg0BJ54cdLa2JX
yk76he1SlG77plz18yf43G8uJW6zRXCHS51tdClom040U9pA0uwiwMf98JtGfdkv7iOjsonnh91K
hlgj3nethNDJWXelIyX4Jz0Vffp8CJfNZKj2bZxT7nRYJkwaE7F1/OC6bA6fqpwKFbZm1EYc2fIn
8Jp5dDRfIGXZAPtJIXcuggE/uFTQOr4g6Jcfm0uOp0rtjKaxegvggkP8hlPEkht7+cb+Pl/VrrtD
ux42Lc2ITIi/ckfySEQ03AeBmHttEdtRvbhL64S/+p2aCp445dppzw4iMubYQuN6O8ahedZKc5t8
OLrY4T+TitaRUWWaZCSrmCH7JzvK1Ssa9x86TVXyHjmfuvM+gmQfFi2cPc3Asny+OO5QUQb8qZ4E
IWhKMpMiFPUypmytui/DDxEQZGGK3PkVPFhw1uI3SsP0B3cNgaQfGDu1O7+xKzYoma/olRxLx0sN
b06C70MBBY1NZlwt3UTSu1vMe8iiDibHpq3U2+uU3F5o1IC0+2CfNem4LsqbSxsu2bmFI/3LtDgU
0KCtAgtNgYq3Dy9LO1y+jpkjbxMktYO8o3LJ7oVV/t+2Z63MbP8yydb3Oh+/00KUJVyqG7mQLgGl
ET6UfP3SxqaNCXJdqNp/LgN0CvJ0H6uMsZiAG1LSUNNr+5Ku/XU5AmD+JoX8Y9p2GJ+LUATH7/AH
NwQbHWIR6ZXvyBIhKA8rICltHoYw5a/RoR6eeRPO6ZBkumPGoP8iS60nWXoD4/HvOi5B3n29bSiA
AwEDTKeSou3/xEW28pkB9CWsxwSLN9935FaQZVQeMYNwi67K92dChXex/+XSq039W7LZdUSjLz1e
mn3ZZbzr2Lsi4xarH+2eTb+YIi3DiZO5ehqWWswWeTIm6+fouMaD52gp+SPU/ALFJKn6LV5hlprB
fX9IlJBydthpMAmHavvPPHxHTpERLn8/xrDXhK56gHVGmzlnweqakN4rBMQsASh9c910h4dWQLAs
6wZXq2kIiJ2sVr/137GhyVfUwxKNZ76obyVIbRPGHFcPoPKF1KMFA5ZDTfavyQiISw6IiZNGR7M/
PQ4DjvRbiEdv0eQOFlOqnNZdA/YLwLPnIL+Nx4n4XInNXy3h7Tkcd3O50H6iYs7mFBDaFo8y0uey
bKalz8k2gIEBKzQyElSZQAstGrx0HCruHfaQujo6cQIOUIA5hcj3/WxBnZy34A8qgnQ0IXhwdFvr
7kcqRxSKmhYpdqXSsJBAMkuRaR/2tFcDHlu1OqUzLk3G6zKcg4BoP7DRPzQdzUNtE5TKN4OoeRsZ
Rva7tPugfdmXfQn/Arrn6NEBmo0kRgtTwTEOAq98LIGsaXLbc1DlkQuD6kVv/bkFOIH3DGcIE6xu
j3qyE0Dx9SX3uWmCrS7N2D3F8WLa4qU8DI2TFzrGmDQy+qyb6qHL36tREP6/Kyco1b7LgB5PJ/aQ
W5zZIScyqdU1JcVQFLW+MKG0SMautb8t8P68tmAjMrYDGQTPOD1sBCCMimW8rJCOt9A5H2Z5enEC
/WeX9uxOdfl3SN+jeuhvl3bF00nPDIUtaFisjl6Uq+erXsYcc7kXvWg4JXuYHsHlQQ/quRbqCnZk
exqHlRGQgE8VCuQZEPoSqQGtO+Y+KM+FaLJH2ubzUBdKkKc4eFI2oLOzxnHFY6SgX61SuAYSFcPO
+HEGf6GORvg+8wpbgWiw4lEaqCyDfyodiyo3ENJzRkDv0F8oULDDD7kLFM/Icq5qiIsoPVtLen3m
DGC3VdTpWB5Ed6GRLg+JGzwyWl5Oc+QGo7Ehtq7VYywQmuONw/QdmLnXl+XXfWDmHtHGbVjAqQ+t
BzRvJ/GTcclrwX6dhtvJvRnisyuQDOm88hn7/OcOmFgj62GzaCMiHZJwggpr2DwXUZuuJp8YkOHm
KwnHsJlfhIl9+POjtSQ3Pyk4aHHhSemQswFyCrsDwGzfjEYbrpvRLu7DEn7wLwSs68AOlEg/+VPM
KQgKcgBJkjEyhzj25DiZXuRLyLCvB0GjI36rgqiu7ZtauZ7RMFekJI2J+knlnRu+n1lX4gtSSoif
AvykA1bEMpVrt804mBtVVsOJoDrcbdE7pcaRxCewSagTX7+UczplPNMNmodXmruniP9TgJEKaQPq
ZbBxEMpADDJfXPxwwbBNE9vS7MENSs0q6oeo39U8b460x4+QKGjGwThHKfXE7O/OQ+YQNtagw5bf
Yk8SJqrnNBNkpprNh6gLjugPFaG/qagjfYCa9BbMVOUCMGPDrRjfnUU2xZhqEwken+dM86m6bp5v
h6DappClqAIBZxM7hD190GW1iwX93PXVXYtU1RLJE5Pl068cisNJaAukH3J9NKkS/4CPfqQoJmcu
I+HAOGcuhqcNBc8u/ie7sw318HOQTIRpAG2EM/73Z006luH3YkIA7Q6s1SaBt1xUEPz6eRuZIe7p
irIGpVqfgXzX19HD7V4XuIyRHmU3zgJZyrD58clDqzdGfB9ZOz4iJYcXgcGTC9dAV4yfBJoMhPt1
G9BmlZOuhRrmo+DV1vUsFhCJgHebyKsPw+IUk+BsV/WIh6XI3Yw1jZchFhYPzyf9s8opfdhx2OaL
PApxe8hUdaRtfOEo/r7CJit3loX/zX1w5Sq+u3QOxsApox6ucLb7khXZVpQ88nQ2KSOPETtG1LtX
QU5wq2Cua7Q0JRvrAwNPWVIwHdkJxPVW0Ac1INN0/RvGzuGFExneCtZDi/vl7rh3Pn2255bzEkr1
haZjjz40wsWlYUCEZUcUDLxfalP2bqfJz3jEDOxHZC/Hb4cGXqHGknurlNLHOL1JJh4TPyTSgQUq
yt7h2/hz3UcrP+1lxRCePwJnGjPli6waYatxIJZ8pdcGUj0nxoUr//JXsAy1S9LpzTqM6zTe0LH+
GyS/GkqqDKufA8ldIX+fAxO/EANsyrCe4zr2D9BwppvYRa3tlM9cx+9UnwOBC32yYGrwXY0HSImH
me0mwT91xbMwygHM8fCFwQAgiU40IEyPuMHEulUhDjvOD4iLx0/eQjbrMS19JR6vad7OjhygG8ot
29U+OpbZNFCp/jjLQCXd0t4tdZl+wnfaGjROZRpfteizFNBPsfYGGsxI88EhM8rVL/HwOst9ZfXm
Nbd6YuFYrDXeYnjRlsnNtllbRcsq1UX9pvz02DK422CaGBUoaHNgFYw+WREMni+5KSBOj3JJshvZ
8Rc+yJ7evPLCqHomnyVbVDt6Dr1fAuq11Kvxkmn503FSXXb7oWPW292KiTZwBXrp6fNgeZAABPP5
P4ueOMxVjdLQOEiCQ7Rp4jv/eLtp4Kj6UB5eKiaaYnMNU6RHz6TrVnW3l81KY0lrAabD49u2WSVe
SFNtrmCiI1cWZF26ydT2K3isX2p8xdrtRAtBOlCAUKTsutRCJw++W+o5Zj/7ho/h6SGtsfJZo8Xm
2159ATf6MAT7H6QgMikZJamdj4cYmE44LYzIqkdPtj/zaG0T0U1KwEZMzqDE9fhQ7EcYmzN+IxKl
EOGFqqBUOQu3lG6vlsrd+/MgzbDpHst+etUSB568t2SYh8LvYgJughGDDid94OYhJGgeG174EWee
KmwpsEl+vohiHIzZiKwB8Yt1NMKcpDiBqlW8YOOrA4JYV2hs+wXZFdEkiKkPrmUkVd3ad0RZ6wKD
OR8VGpvCuBFVh7suHCj95sRe7wbHZZ5vYsYYOPfo1KH0ttxurnz0LARlTWTeMXIzra/6NWAShM8R
ZC73kFjYKk49Ua2KBdSiYFvikE/y06NXlOla37Gsi2PlS/sYPwKZVzoxOuOFhfUz1eV+bKIhtH3N
OuzMA2hUW+kNr6wpdehXzcpYVPq6CYg9L3HQDxjhK2lLdcQpWGc/O4mvb3+PXrLU6+gjcOvjbxwe
xFMyDkNLOkaoLtb5B0bbSKiQD0Mcosry27H+5aLpkFMrOzW+xisLKqRuKOQgOAbk0wjgknO5/psG
jWWyCi6eJOWSYNjyydLVxeHc3Wxtxu0zPX6cA+qSUTTCpWcn6BE7RMANmLoDd4bxrRtxjNuuEVPk
6Rjf5eeg3dHmNoPggc6UayYpLXt+gCswnOZTkNms0DatFAIyq1vkC1laMTYsJXij1LfuPVIwK3SX
Z9z2nWg/ecCz/Z3+bq/0Ya0+X6e0J7PN42glxBtLGgzSSSVirgp6L08pvnJfZiAU61ArjiIHlZeP
AFHA/I5eZbLdAd9TNSkw9H0jj7yYuNLjhzKqiQcxjdT17M7O1CDDC4IWuA2hpzuCqfd5NUdKytCm
/iddWU1K8bBdsVjmeyZJ/fDRm7wQEq8DJlHcT+BrVR/2p4Sn/yjeJZH9CIRiMLzn5KI98qgStKkT
Qj0mVieOvcyZimOH7HcVxV9lP9407AHx8TV8gake4UrDaJmXJZJEaco/8SsORqEuzWV6Vak4feZL
k1gDvuaCmXYUqcwjdJB4Ai82bPdbUzSVFAOxOKEGfAH8wm8U6lu+j+W7MHz3frtqZf4pxXSeZ0CI
8SccyRnB61Rrq770b4O1Cp8Fcx8ON5ZEmod8ZrMePKy3Jt9s/T+YoLl4nZL5JaWKoGLOnDByRWwk
foy155jzQDN+YzQE77vMOUTc8ogP+VN77codgArwDlJmSS1m8EV7XdNUVncmOURQd3pOxy/U5kug
0ZUr4xJhuOPp0Y8O3BOKaGnYrqQguK1yo1GgOiMi6n5N6LIJYMgQu7C4R4pSaCSRQm2W6LiNN7WP
LWZpWV+NYkhtGWEfi5xFf3O4LAVhLU4mDWFlUc+1u3ckIOW53xgE1mPODqM4DuS3Rpy7VjCRZNhb
XWk+/lMaZDdL99od4WVefcPgrDacEQqwHPDpYZJEY5KJOeBZXFDuSKjFTnlOYgf7ElN5L0Qsu8i4
d/2YAcxayTTVTXPG4zm1qfZAgENALMvyuGNm6eRE14voi7jd2DGBihwkWJN8oRAI8TwNau/7g5gM
ckHPcn0swnYXUwqkh1EcOQerZVxINpKO05Pf4ZkhBP9h8I80DveIIaHzUH220dw6vXCLJAvnRu4c
1ZaVwcWcpixQnwlKOWvswNzqkkcsXV43x1PsR0DmlyxHq6UQrejlyZb3o5QFqATbCYEBDuNLEmws
YIkTNd8noprDWkiWRqlnqOPNubTDyhPhbRreWcLRmVSVXC+eGU5Us/yWywB2htpODbd/5gSmHM02
XeW8gLQsqCsSyngMmRtYwciS5B0Ur44e55ARfYiQ1ImyTeaAY2ukVQI5D1H3iS9Nw8apBUjm8nuf
UTWibLGDgfkb8ENlw0Y5+gXePNv8VcNBJzGDPYbi2Ii+isgUKJO6DoVzVPIHQES0R+S7xCK/mT4G
W7KaEEizKrP2oANg4Orp/1iP+hmqZF4VdHrFDHbJ8A5MMsfv34cMiHpFFXHSpzFv4gr2ck9w4KrT
OiD5dyO1CXhfP968U0XzpB+huXyTBurK6o5FRyEZH+OtgxnuE6GKHskSFC970+roTG6sg6Q/4xif
vTIubnz7POGk7dTJgHspdgryPt950JGm21B1zTMgw2EhQox/n/xmSFCtEXYjJqURkWikfXkNHnKO
avJHHTSdATzhu9aUNWWIEdz6wJgwL1wfg/6vMDzqlSgLRfjrjMyQkWAIqJrefn+K3kly2JbCyzSV
o6N0AxlUXb8XXpessPAhConmwUoDjnzkpS1OTbQackYIqLYbLhhHXaufCJAQdmlZE8pLwOJnzRHA
4UEBN3eItvRJ5wFc8ZcAA2/0u32KBb23ayyBaLlko/fmC6BTJx6vuG5mcM3Olw5wrN7Mvwpo0MVi
113jdpIFCAit6epUMYJkehaODYp94TbJKzzmaeK7ytCuWtR1TLVyy/dHsaKwkE799CIaaak7MUuT
d7YBSJn7zqgW5KnZp29sIYBUvzoqjyrHYH0TERiy5+1u0VfHWc2NMhIiMyCKTloshLHh22ZjNtsD
dSJHLoo3ADaXICNWW7LKSWUAHuS7dndoCaTcjdY9zZUwAjpW1qIK6NYbN29pFezX4iYtWz9XB9v4
ijYlWyVY1pXmu2PlRm/Fj4skaJmp7Z0pdvhf+sOrp+j+afhQwQjOJawGiABvtcltZ0bxRfqsTLcc
2p5c03Zj4RsE3jLQ4SMWIwzuGU/IHOpFcKmJq9dl3y9WTB8FcoM5idvNL2b1AvxAcM3zeOC8w7yu
qcpIkS3593PaLXU0IRCl5o2HAJ2hWWJ35uk1ykyX3ptnyEbKRN28KJlnCUW59dNiekb9VYymau0e
pCE6OwftEHnojPGGjAWkQLXWB2rDNUUFvf20lJ5IcUCfrHfPkE9NqFut4FM5UfJXQQFmioVd1BRy
6S6VmkQs7S1sJD16xtj5TTMeaAoQRn663hSS9HKKDFsac0jvGTmmOxlMt6Xdoxj1eqZ4CRifkabU
KaqfHNH+O6KO8H4zLv+6KyXHBi7OwUrdPXbzAl8yME/yaOy20pia1UvfmYhjfD3U+RitGDuE+3sq
kXXn8oaB9M1mFVayTExHUa0z2UXETiltyYget/Mrb3EtsE4KZ0HRm6/JEFhx2WMcuh3bTqvdeadx
X2MVBG5nR+K+Ri8tDOVHL6FIucXO4z90r6Va9XRw4u/xYl+9Hrz/muI03/IYFTlnprzV4fvOZNQs
wOP17VvBsjoF8OI9ktRdxR9kuqWKRXBQnRNsfW/dbDKPxNzpJR5030iU90GGGzSursMYOfXBxZMi
Ibe4cUQBlBiyXfLmo+p98OvSB8cCSfL0uxWydg0AAw533zAAtQG946N/M4h5xJ50MMQgARCXGnb0
vrLk7q55vwe4eYneVMWmAVZoy9KFOC52JmVIRrsN7KWXur2vDQEtdAUUN2LTKUo9Er3er5DkcolX
Yr/QlJDUjquzujCeiz3oVm0fL0JGokf4+caUFcG+2/B0oxhQZnokhuSON5Sph3Xy40/MvSFatcHh
oTFEr3J4VQLTV1qE5MAHFdzfmGKKTjn8iw5w+7Fvv9UzC7QJ3SeqKeTx5jOkr/fu7vMI6Ji2jdQE
U5Q0UzYZE2NqKDp4sKTyVbe3Xr+IReykRndqnT92Q5PkIsjjQqIavcoQM4SQQBWFZav6vtpx0cI2
hs7V8Dd7wqN/+Ka9XN8ucuIFpdxlxhKjASKxQb+Q+r6etMrzQ3pydF1aeKHtLMmm5jFNH4zd9VLr
bHUcPQWj/yMrZKo3sN0SQB/vK653CvOEBuwM43PxBRPrhAievpT7PQ1gJqIMkdqE1DQavo0Cjsvx
Z5odQKRrsTle0IJUAKEGf5KcWALl5kc5SKJxBjkQbdrb6aQwt2cUPDlXaRKhLqztU3E0zZtD1BSX
mIfAMOwLXIztIogKNwjADrGe6whmQFKMdXs1RWjeX502kk2Zo/LO8ZpARw4wrKVjy8yQA7D1wN+O
U2Ula+0zNELJJg1plceMbPQ9LrrPYI61lVwFHDqGpAbk+++1elklnoeh3W/sQcNNiAHnzEl1KN3O
2U/L3YBJQduiDVUaZ1KvNCmPF1+DQQnM0plUXcekeGnma4yyBgKuKeCemtY5Zg0e0TpFTlaZBnCw
AaLw78OIXjsG80FAgFNjdXULiEvWsmdYqpMq7KZMMWD3vd8XozgLyNuGb+yE9u8Kv6slc/AJD+Dg
bEgr0vt+VqoXXJ9U64Xpj2TDGb7muDqxzUh8jRMsd4wHGfA+rg6cce+AuK3hTNyEr2nAIIGzIK/H
W7Xxt2sCo5kjShEv5bp1eU1RyiXFju8qFrtwDSEMmlSwofp06f6s8nfRpmG6cWDdRxma+o5v0FhN
SJQSqUMsU/S/kqHsRBOJeMquwxOGJ3XcGM+Kud73SmrHEm5XlZSzQYRbvEfc5/rx2aR44CD3ZPeM
OGCC+lbGEIISezXNTZiLZD8XvN/jzrMuOCuvX3NlWhQhBTIKx5PwU2yxvfvleoMdRmVTnVVe5xcq
UM/YJSnlKI+/SuPBP1f236bBILmpb1cd9WaWAYW0H4fC7b1zcafQnbSfeZszqg4pGMbdNMlE9DsS
D0rFwHpSe7DSop09n8w5ENJXtQW/bsdv3OoWZpnJKoEU9ii0qBCcXH2V1naSmnfR2o7qXfmIgeae
fcKCi5O/vGF6cCoXMQFjYBTkdFOk8Ycttivet/DS47+2KcvDcD1aLl5nKEWW2b3iv8qbXYaJ8q+b
sJM4ckQnpt5OtBM/gsdIZpDM34D0Os5py0fcHGtgWbsLczU4DM3smfbKJLo1/vHCoUiVU87dsabp
TMKqNu+UoWDvQJaChgnUGLI6kAzqA3Y/1HXjNg58+uVtXb3lhtPCLriPPzD51vMz2VOq+zrMU3tA
nddIeRw/nguvzqw8PHu+F4oGJK/hGRjMigxKkI223gQ55U0HPoYN2Xnu4BRIQcc0LemvN1q8GZ5y
QSsWAR5NJ5wz7GJuFq/Wfzelsw8qOaeWMiXpPd1k3U9fFLTio3BB88rocmjoqvOVIV2aoMIDLzcH
1o/8S6evJa3dDCVBqkZJpWWHRB2Yvj4R7WTRdQFL7TawXxpK2WRknwinm02HNv5Ctjan5MlcMs9+
W8k7cuDHfN+7zr4xnlp4lD2TcC/n1tJb5uApH8w/B4qfZfDTbH27IvIjzIY3Kp/LWvn8ixrtxFS4
lv7Hn8yYR3LKoTntkpdmBlSZhyCt04WjlWnRN6Sq3/2aY5FyyUUQ+zTPW0ksuNoUwgVhL5fxIHYU
5I3XHkCuL7H4Xa0daAiOeKWoeBsh6CZvdHu6Yvgg9k9spWzIYkiYsBgq5SlBiCF6Ne+3V7bnAc5J
vpaLR79om4DGXDioE4YkhZCfkeCKOgK6v2xOAQXSh3PEhHYxVHIkZXrGnyScdn49LZlqeDeTleXg
vAkEEFdwdnx63lJ+DAHElgtPT+cvM7yErWY5w93CLA2RiYEMJ8pjTnLaNDWT6f3gf4byK8o9WS9m
W857NMhzHkkT+3OA88mEx4InLoRV69c19kSV+MAsynbHnPLzZry8CewNyhV/DY1hDa3IZiQERrDB
zx8mr84o0qdrU4eBaLW9wTZf2nYd4bb3hRFsfQl9yR+YJ6d6usHoZS9BnRNQZjqXuOcvsHstfeel
BsujiS3y0PXPogirTlHZKVJi8yxVmrOM73Npc1YeyX8rRcGR5qy5+t+noZwEqw/H0lJYfUuj1Fu9
ud70DnlO/ZJtXfN3YzJ0x5MpKS1vHxIRAQNTzcXwbXnlVXSoU4A3N91j5f3zQcjc3oD4d4Rml1Xa
G3II8C42/OKD+LRxmEH7bRvLA2G0CjS1azkd2XtNIi0tbMhgMMa6NDNTXBuqv3aBqZm0flSMc0Mj
+9tVlKcKH5QVBn2vjahPQmwm58sCLZbOtaZ4fFdmxkZ5mVekdjhHHV1+m2R4US+/G3WF9FEAeyO0
BnEZ17JEjrKWj3pHhqJonU1PcxveL7dA8mdrNYMEwZ263ostijXX6G28lpOWQ9WDLVofDSdta/HX
ws2yyK68lE2YJpua8M0IXSrMPU+r1k3rLdUJJLRTedwIRhLx2XCo4x7G8T/U8AE4HIFBaDoPEZFa
41m7NlwviJzJ97rs3p6hjJLB3M9QRdFYnl/zJe5W0AY7cnvYgdA3knbm9PmcmVEuLDS7S7/gJu9M
+BdtACrWhLPhimtq/1i5oOIUVYoT6e3DrYJA/qdS8Sa9kwnrQl9kfhgD7XRqkdJmiKggxfqy3aHd
UwCjPDbQ9jCf40p4adj3MgRw4hhPhNHKof5ke1dMPP4eeNKn/wpkWnhoBP7KSmTfBZLy6f55mTro
Pk7fBys9sKSVgcaoTdq8APhlbSvPpFDuKioFGDhmdXsSOrvy9Z8PIF7Qv4pGZMWfXnpH/O9iyx/T
W3r94rjaBC9ZYj2DMU0lLU+ap0Oj8blFZg45WnU8qtzq72tgPxg3zb04EDPViaRM6LWGuLuFg27B
uoojQoLi1aEre4VGREqT3yaqxrMvWbxpyVobLm0h1nazazXgWq4gHGl6eggjUvZoGSSub/0fmlf+
0xaO3oI0Zz8YvMEURSsxoYy4f/7jFRoEfTdL72iKRAP5M0q9FCdkRJtsHAlT4WkIR1/rZDD37GHw
4/SZwRtelaXhmX3GwG7DmCKAtUTYVGIiBstA/qrK6yziCwrz63xLJnlNnJ+ffnpFrX8KU2m9cYds
JQp/RM3Gvhl1xIOoDksjcIYT4uDgK+cAJlT39V7+0WKhm0/X6XDwKqWa9K/I+d5MFhMN5pC+xiVh
1Oyyqt87ypIZvHYwPuZrZ3KohGNnxL5L8AK3pYHYr29GCr/KrTSUzR+a5r/IRN1K3wnz9x+c5/Gj
26JB9zLU7+bBLAl1LJFUd5xfVVpJANekqpfbVOc4boW+f000rnzOf4GrEsQYeJRJzjIscjfvCl7W
AcCWrms0iGTHuMitXD1LoVggHxOANoB921We16a9bpVBMZrGCAaYjDri2k25oSojvJ2nRPCU9QgN
y3NMXG+Hf+/Ek9KntfM8FvGFqQ3NY74hfqNGoPE5M8Qmwem7MBGqUn0vimqQ5moUoofZjAgUylEZ
FRjzfg4fwowyZdCKoFbLka7Ezfye0P0IyksIp9d428cfP0NGqyA/xoeRXR90Q+Cbi5DFmcvbkADj
kzepFdX6Give+C+Ej2re2rguxkH2S5HrL5lNPRr/g+XAHARqGPF3Gx/MOpQmou6sKREBAdBCmJGZ
c1naGCgMKFG4XgmY5NkjkdDV+9QMyvZNRyQ5UA4ovszdk8uYfwUsFB9p9TKQfw7b7ihrIE0/AoBf
ORLxGhjo28enkHFq/AA3QaWupkIj/lXij4Y2gtFKz5+VmULOoEJXQBZpd9U1lRhWV7b6yq5v9EPM
/EnbtYZSuhVF68rJYjUEHanziVhk9XkBOb4fuRgRa/gvX9qIDuhPckMGLa4UzW1ggD9mBOVb/VyO
7ZGWiYTOFlaWstn0FlUUs9JL6knIX4kmKqp1eIjiO8JCIm5AFtQilGmCSqNOrz2PPdH6PFzGif7C
ZFV+WO25BhQoQWzWHhsa8TGeKbXs1tXTXMt++X4pMI2Y0eCr3mLXZ4ic2T1LNnh6+/140NFTrO+8
/zpvIkBoz2+8mW6huY7W/i/1R+lPf9wsxAGp5tLTJ00gxLgoqV7Obx+o3qwHpT7QPyFcp2ImJsdh
KDrb4xEMI2ejrDBQZ7v4wpl6pSveCtVO4ierX//f0PKmYzQbsrulHa2FKri0UwRwHfDjGknWQZmM
shGsAPefrMmgirDvIq5NwJrNTXvOelKFqz3bJRyN1pquKrI0+atVIzks46irWgOlWQCQNelZfAm+
WozBhaQrFFnSvuLMcM55XcaJ/TFweuZeLwvvvY4vw5Dh04nvYNaNQSq/X4jPVFDXbl3J/feJA+60
YR4TuZXLPCd3nnwZtfWn71ryVo8QzcezO5GXhO+VyqrJPLCb54v8EbLGBvyOLN6H96xGu6xa503T
US6Iql9QKbBcIERtFGUZhRXf0mDJP6zpNEKU9G+0wzsyhDZXshCbzBhDp8bSJDXTNqoIovhrxaAn
DStgaiG0MIh62XXiK9sXzofiPmDSXApQi8VKasMqmSXrTW/nvLSX7moJqLKFfK4kyTfCAJwIcooj
FXRoVcVS4tLBNRq1A9WIqvy4A8Eiq7tT8WvNM+vH9hflx9h4GcKHNkZqhDM5xGV6vh8pZJICOwES
Nv5tYbNLzt15r3xPEG89v6BvEWcDqf1SuLQW97Cwb+A6IaQELleJt8Flo2koADmcMZJ1R4XvFZAK
IXEougfw
`pragma protect end_protected

